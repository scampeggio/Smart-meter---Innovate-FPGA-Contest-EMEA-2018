library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.std_logic_signed.all;
use ieee.numeric_std.all;

entity vga_generator1 is
port
( clk: in std_logic;                
  reset_n: in std_logic;

  STATUS: 	in std_logic_vector(15 downto 0);
  FORCED: 	in std_logic_vector(15 downto 0);
  CHARGE: 	in std_logic_vector(7 downto 0);
  DISCHARGE: in std_logic_vector(7 downto 0);
  P_SOURCED: in std_logic_vector(7 downto 0);
  P_SINKED:	in std_logic_vector(7 downto 0);
  BATTERY:	in std_logic_vector(7 downto 0);	
  
  h_total: in std_logic_vector(11 downto 0);           
  h_sync: in std_logic_vector(11 downto 0);           
  h_start: in std_logic_vector(11 downto 0);             
  h_end : in std_logic_vector(11 downto 0);                                                  
  v_total: in std_logic_vector(11 downto 0);           
  v_sync: in std_logic_vector(11 downto 0);            
  v_start: in std_logic_vector(11 downto 0);           
  v_end: in std_logic_vector(11 downto 0); 
  v_active_14: in std_logic_vector(11 downto 0); 
  v_active_24: in std_logic_vector(11 downto 0); 
  v_active_34: in std_logic_vector(11 downto 0); 
  vga_hs: out std_logic;             
  vga_vs: out std_logic;            
  vga_de: out std_logic; 
  vga_r: out std_logic_vector(7 downto 0); 
  vga_g: out std_logic_vector(7 downto 0);
  vga_b: out std_logic_vector(7 downto 0)  
);
end vga_generator1;

architecture BEH of vga_generator1 is


-- Images
type LOGO is array (0 to 119) of std_logic_vector (0 to 249);
constant GIORGI: LOGO:= (
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111100111111110001111110001111111111111111111011111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111110011111111001111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111000011111100011111100011111111111111111110001111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111100001111110001111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111000111111000111111000111111111111111111100001111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111100011111100011111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111000110000000000000000011111111111111111100011111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111100011000000001111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111100011111111111111111111111111011111111111111100111111111111111111111111111111110001111111111111111111111111111111111111111111111110000000001111111",
"1111111110001110111111111100001110111111111100001111111111111111111111111110111000000000000000000111110000011111111001111111000011110011000111111100000111111111011111111111111111111000001111111100001111111111111111111111111111111011110000000011111111",
"1111111100001100011000111000001100011001111000001100111001111111111111111000011000000000000000000111100000011111100001111100000011100000000011111000000111111100011111111111111111100000011111110000001111100001100011111111111111100001100000000011111111",
"1111111000001000010000111000011000110001111000011000110001111111111111110000111111000111111000111110000001100111100001111000000001000000000011100000011001111000011111111111111111000001100011100000000111000011000011111111111111000011111100011111111111",
"1111110000011000110000110000010000100001110000110000100001111111111111100000111110001111110001111100000111000111000011110000000001000000000111000001110001110000011111111111111110000011000011000000000111000011000111111111111110000011111000111111111111",
"1111110000110000100001100000110001100001100000100001100001111111111111100001111100011111100011111000001110000110000011100000100001000010001110000011100001100000111111111111111100001110000111000010000110000110000111111111111110000111110001111111111111",
"1111100001100001100001100001100001100011000001100001000011111111111111000011111000011111000011111000011100001110000111100011100011100110001110000111000001100001111111111111111000011100000110000110000100001110001111111111111100001111100001111111111111",
"1111000011000001100011000011000001000011000011000011000011111111111111000111110000111110000011110000111000001100001111000011000011001100011100001110000011000011111111111111111000111100001110001110001100011100001111111111111100011111000011111111111111",
"1111000110000011000000000110000011000000000110000011000000111111111111000111100000111100000111100001110000011000011111000111000010011100111100011100000011000111110111111111111000110000001100001100001000011100001011111111111100011110000011110011111111",
"1111000100000011000000000100000010000000000100000010000000111001111111000111000000111000000111000001100000010000011100000111000000111000110000011000000100000011000111001111111001100000011000011110000000011000000011100111111100011100000011100111111111",
"1111000000000000001011000000000000011011000000000000010011110001111111000000001000000011000000010000000100000100000000000010000011111000000100000001000001000000001110001111111000000000000010001000000100000001011111000111111100000000100000001111111111",
"1111100000100000011111000000100000111111000000100000111111110001111111000000010000000110000000111000001100001110000001100000001111111000001110000011000011100000011110001111111000000100001110000000111100000011111111000111111100000001000000011111111111",
"1111100001100000111111100001100001111111100001100001111111100011111111100000110000001110000001111000011000011110000011110000011111111000011111000110000111100000111100011111111100011100011111000001111110000111111111001111111110000011000000111111111111",
"1111111111110011111111110111110011111111110111110111111111110111111111110011111000111111000111111111110001111111001111111111111111111111111111111100011111110011111110111111111111111000111111111111111111001111111111011111111111001111100011111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111000011111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111110000111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111111100001111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111000001111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111000011111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111110000111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111001111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111000000000000000001000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111100000000000000000011000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111110000000000000000001111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111100000000000000000000111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111000000000000000000000111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111110000000000000000000000111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111000001100000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111110000001110000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111100000111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111100000111111000000000011111111110000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111000000011111000000011111111111111110000000000001000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111110000000011111000001111111111111111111100000000011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111110000000010011000011111111111111111111111000000011100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111100000000000000000111111100000000000011111100000011100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111100000000000000001111110000000000000000011100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111000000000000000011111000000000000000000011110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111000000000000000111110000001111111111100111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111110000000000000001111100000011111111111111111111100000000000000111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111110111111111011111111111111110000001111111111111111111111111111",
"1111111111111111111111111111111111110000000000000001111000000111111111111111111111110000000000000111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111",
"1111111111111111111111111111111111110000000000000011111000001111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111111111111111111111111",
"1111111111111111111111111111111111110000000000000011110000011111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111100000111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111100000111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111100001111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111101111111111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111100000000000001111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111100000010000001111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111000000111000001111000011111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111100111111111111110000000000000111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111000001111000001111000011111111111111111111111111111111111111111111111000000011111111111110000000000000000011111111111111111111111100000000111111111111000000000000000001111111111111110000000111111111111111111111111111",
"1111111111111111111111111111111111000111111111001110000011111111111110000000000000000000000000000111111000000001111111111000000000000000000001111111111111111111100000000000111111111100000000000000000000011111111111110000000011111111111111111111111111",
"1111111111111111111111111111111111000011111110001110000011111111111110000000000000000000000000000111111000000000111111110000000000000000000000111111111111111111000000000000111111111000000000000000000000000111111111110000000001111111111111111111111111",
"1111111111111111111111111111111111000001111100001110000011111111111110000000000000000000000000000111111000000000111111100000000000000000000000011111111111111100000000000000111111110000000000000000000000000011111111110000000001111111111111111111111111",
"1111111111111111111111111111111111000001111100001111000011111111111110000000000000000000000000000111111000000000111111100000000000000000000000001111111111111000000000000000111111110000000000000000000000000001111111110000000001111111111111111111111111",
"1111111111111111111111111111111111000001111100001111000011111111111110000000000000000000000000000111111000000000111111000000000000000000000000000111111111110000000000000000111111100000000000000000000000000001111111110000000001111111111111111111111111",
"1111111111111111111111111111111111000001000100001111000011111111111110000000000000000000000000000111111000000000111110000000000001111100000000000111111111110000000000000000111111000000000000111111000000000000111111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000001111000001111111111111000000000000000000000000000111111000000000111110000000000111111111000000000011111111100000000000000000111111000000000011111111100000000000111111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111000001111111111111000000000000000000000000000111111000000000111110000000001111111111100000000011111111000000000000011111111111000000000111111111110000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111000001111111111111100000000000000000000000000111111000000000111100000000011111111111100000000001111111000000000001111111111111000000000111111111111000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111100001111111111111111000000000000000000000000111111000000000111100000000011111111111110000000001111111000000000011111111111110000000001111111111111000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111100000111111111111111000001111110000000000000111111000000000111100000000011111111111110000000001111110000000000111111111111110000000001111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111100000000000000111100000111111111111111000001111110000000000000111111000000000111100000000111111111111110000000001111110000000001111111111111110000000001111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111110000000000000011110000011111111111111000001111110000000000000111111000000000111100000000111111111111111000000000111110000000001111111111111110000000011111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111110000000000000011110000001111111111111000001111110000000000000111111000000000111000000000111111111111111000000000111110000000001111111111111110000000011111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111110000000000000001111000000111111111111000001111100000000000000111111000000000111000000000111111111111111000000000111110000000001111111111111110000000011111111111111110000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111000000000000001111100000001111111111000001111100000000000000111111000000000111000000000111111111111111000000000111110000000001111111111111110000000011111111111111110000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111000000000000000111110000000001110000000001111000001100000000111111000000000111000000000111111111111111000000000111110000000001111111111111110000000011111111111111110000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111000000000000000011111000000000000000000001110000011110000000111111000000000111000000000111111111111111000000000111110000000001111111111111110000000011111111111111110000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111100000000000000001111110000000000000000011110000011100000000111111000000000111100000000111111111111111000000000111110000000001111111111111110000000011111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111100000000000000000111111110000000000111111100000011100000000111111000000000111100000000111111111111110000000001111110000000001111111111111110000000011111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111110000000001100000011111111111111111111111000000000000000000111111000000000111100000000111111111111110000000001111110000000001111111111111110000000011111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111110000000011110000001111111111111111111100000000000000000000111111000000000111100000000011111111111110000000001111110000000001111111111111110000000001111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111000000111111100000011111111111111110000000000000000000000111111000000000111100000000011111111111110000000001111110000000001111111111111110000000001111111111111100000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111100000111111000000000001111111110000000000000000000000000111111000000000111100000000001111111111100000000001111110000000001111111111111111000000001111111111111000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111110000011111000000000000000000000000000000000000000000000111111000000000111110000000001111111111000000000011111110000000001111111111111111000000000111111111110000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111110000011111000000000000000000000000000000000000000000000111111000000000111110000000000111111110000000000011111110000000001111111111111111000000000011111111100000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111111000000000000000000000000001000000000000000000000000000111111000000000111111000000000001111000000000000111111110000000001111111111111111100000000000011110000000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111111100000000000000000000000011000000000000000100000000000111111000000000111111000000000000000000000000000111111110000000001111111111111111100000000000000000000000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111111111000000000000000000001111110000000000001110000000000111111000000000111111100000000000000000000000001111111110000000001111111111111111110000000000000000000000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111111111100000000000000000000111100000000000011110000000000111111000000000111111100000000000000000000000011111111110000000001111111111111111111000000000000000000000000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111111111110000000000000000000111100000000000111110000000000111111000000000111111110000000000000000000000111111111110000000001111111111111111111100000000000000000110000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111111111111100000000000000000110100000000011111111000000000111111000000000111111111100000000000000000001111111111110000000001111111111111111111110000000000000000110000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111111111111111000000000000000000000000001111111111100000000111111000000000111111111111000000000000000111111111111110000000001111111111111111111111100000000000011110000000011111110000000001111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111000000001111100000000011111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111000000000011111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111110000000000011111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
"1111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
"1111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111000000000000000011111111111111111111111111111111111111111111111100000000000000011111111111110000000000000000000000000000000000001111111111111111111111111111111",
"1111111111111111111111111111111111111111100000000000000000000000000011111111111111111111111111111000000000000111111111111111111111111111111111111111111100000000000011111111111111111111110000000000000000000000000000000000111111111111111111111111111111",
"1111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111111100000000001111111111111111111111111111111111111110000000000111111111111111111111111111111000011100000000000000000000000001111111111111111111111111111",
"1111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111110000000011111111111111111111111111111111111000000001111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111",
"1111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111110000000011111111111111111111111111111100000001111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111",
"1111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111000000111111111111111111111111100000011111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111",
"1111111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111000001111111111111111111110000011111111111111111111111111111111111111111111111111111111111100000000000000001111111111111111111111111111",
"1111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111100001111111111111110000111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111111111",
"1111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111110011111111111001111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111111111111111111111111",
"1111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111"
);

type IMAGES is array (0 to 14) of std_logic_vector(0 to 151);
type SH_IMAGES is array (0 to 14) of std_logic_vector(0 to 79);

constant AVAIL: IMAGES := (x"00000000000000000000000000000000000000",
									x"00000000000000000000000000000000000000",
									x"03e0e0383e03f8e0003fe01f01c1c38ffc7fc0",
									x"03e0f0783e03f8e0003ff07fc1c3c38ffc7fe0",
									x"03e070703f03f8e0003ff8ffe0e3e38ff87ff0",
									x"07f070707f00e0e0003839e0f0e3e38e0078f0",
									x"077038f07700e0e0003839c070e3e70f0078f0",
									x"0f7838e0f380e0e0003c79c07867670ff87fe0",
									x"0e383ce0e380e0e0003ff1c07876770ff87fc0",
									x"0e381dc0e3c0e0e0003fe1c07076770f007fc0",
									x"1ffc1fc1ffc0e0e0003c01e0707e3e0e0079e0",
									x"1ffc0f81ffc0f0e0003800f1f03e3e0f0078e0",
									x"3c1e0f83c1e3f8ff8038007fe03c3e0ffc78f0",
									x"380e0f8380e3f8ff8038003f803c1c0ffc7878",
									x"00000000000000000000000000000000000000");
									
constant USED: IMAGES := (x"00000000000000000000000000000000000000",
									x"381c0301ff87f00007f000e00e0e063ff07f00",
									x"381c3ff1ff87fe0007fe07fc0e0f0e3ff8ffe0",
									x"381c7ff1ff8fff8007ff0ffe0f0f0e3ff8ffe0",
									x"381c7031e00f03c007071e0f071f0e3c00f0f0",
									x"381c7801e00701c007079c07871f1c3c00f0f0",
									x"381c7f81ff8701e007073c07871b9c3ff0f9e0",
									x"381c3fe1ff8701e007ff3c0383bb9c3ff0ffc0",
									x"381c07f1e00701e007fe3c0783b99c3c00ff80",
									x"381c0079e00701c007f01c0783f1f83c00f3c0",
									x"3c3c4071e00703c007001e0f03f1f83c00f1e0",
									x"3ff87ff1ff87ff8007000ffe01f0f83ff8f0f0",
									x"1ff07fe1ff87fe00070007fc01e0f03ff8f0f8",
									x"01800e01ff87f000070000e001e0703ff07038",
									x"00000000000000000000000000000000000000");
									
constant BATCHARGE: IMAGES := (x"00000000000000000000000000000000000000",
										x"00000000000000000000000000000000000000",
										x"3f81c3fe01f3870707e03e1f3860fc03f0c718",
										x"3f83c3fe03fb870707f07f1f3c61fe03f8c718",
										x"31c3c070071b870f8770f18e3c63c6031cc718",
										x"31c3e0700e03870f8630c00e3e6300031ce738",
										x"318760700e03ff0d8631c00e376300031cefb0",
										x"3f8660700e03ff1dc7f1c00e37670003b86db0",
										x"3fc670700e03ff18c7e1cf8e33e73e03f86db0",
										x"30cff0700e03871fc7e0cf8e31e33e03e07df0",
										x"30cff070060b873fe670e38e31e38e030078e0",
										x"3fcff07007fb873fe638ff9f30e1fe030038e0",
										x"3f9c387003fb873066387f1f30e1fe030038e0",
										x"3e18186000c1873066181c1f306030030030e0",
										x"00000000000000000000000000000000000000");
								
constant BATDISCHARGE: IMAGES := (x"00000000000000000000000000000000000000",
											x"7c0c3f81c0f0402184183c030f1840803c3108",
											x"7e0e3f83f8f9f0f98e1c3e0fcf9843e07e3198",
											x"7f0e3f83f8f9f9f98e1c3f0fcf9c47f07f3398",
											x"631e06031c6309898e3c331c471c4e10733398",
											x"631e06030c6303018e3c3318061e4c00731398",
											x"661b06030c63c301fe36331806164c00731398",
											x"7e1306030e61f301fe363f3806174c00771ad0",
											x"7f3306030e60fb01fe663e3bc613ccf07f1af0",
											x"633b06030c603b018e763e1bc613ccf07e1ef0",
											x"633f06030c601b818e7f3618c611cc70701e70",
											x"673f86039c7339c98e7f331cc711c770700e70",
											x"7f718603f8fbf1f98ee3330fcf90c7f0700c70",
											x"7e618603f0f9e0f98ec33387cf90c3e0700c60",
											x"00000000000000000000000000000000000000");	
											
constant BATSTATUS: IMAGES := (x"00000000000000000000000000000000000000",
										x"3e00e0ffbff7f8f81c3800c1ff0607fce1c0c0",
										x"7fc0e0fffff7f8fe1c3803f3ff0f0ffce1c3f8",
										x"7fc1f0fffff7f8ff0e7007fbff0f0ffce1c7f8",
										x"71c1f01c038700e70e700e18380f80e0e1ce18",
										x"70c1f01c038700c707e00e00381f80e0e1ce00",
										x"71c3b81c0387f8e707e00f80381980e0e1c780",
										x"7f83381c0387f8fe03c007f03819c0e0e1c7f0",
										x"7fc3381c0387f8fe03c003f83839c0e0e1c3f8",
										x"70e7bc1c038700fe01c000783839c0e0e1c038",
										x"70e7fc1c038700ce01c00038383fc0e0e1c018",
										x"71e7fc1c038700c701c00e38387fe0e0f38e38",
										x"7fce0c1c0387f8c781c00ff03870e0e07f8ff8",
										x"7f8e0e1c0387f8c381c007e0386060e03f07e0",
										x"00000000000000000000000000000000000000");
										
constant LOADS: SH_IMAGES := (x"00000000000000000000",
										x"00000000000000000000",
										x"3c001fc007c07fe007f0",
										x"3c007ff00fc07ff81ffc",
										x"3c00f8780fc0787c3c1c",
										x"3c00e03c1fe0781e3c00",
										x"3c01e01c1ee0780e3f00",
										x"3c01e01e3cf0780f1ff8",
										x"3c01e01c3c70780e07fc",
										x"3c01e01c3ff8781e003c",
										x"3c00f03c7ff8783e203c",
										x"3ff87ff87ffc7ffc3ffc",
										x"3ff83ff0f03c7ff03ff8",
										x"1ff80700e01c7f000380",
										x"00000000000000000000");
										

--//=======================================================
--//  Signal declarations
--//=======================================================
signal h_count: std_logic_vector(11 downto 0);
signal pixel_x: std_logic_vector(7 downto 0);
signal v_count: std_logic_vector(11 downto 0);
signal h_act: std_logic; 
signal h_act_d: std_logic;
signal v_act,v_act_d,pre_vga_de,h_max, hs_end, hr_start, hr_end,v_max, vs_end, vr_start, vr_end,
		 v_act_14, v_act_24, v_act_34,boarder: std_logic;
SIGNAL color_mode: std_logic_vector(3 downto 0);
signal H_CNT,V_CNT,V_ST,H_ST,V_EN,H_EN: integer range 0 to 4095;
signal PHASE: natural range 0 to 10000000;
signal PHASE_CNT: std_logic_vector (7 downto 0);

begin -- BEH


H_CNT	<= to_integer(unsigned(h_count));
V_CNT <= to_integer(unsigned(v_count));
H_ST	<= to_integer(unsigned(h_start));
V_ST	<= to_integer(unsigned(V_start));
H_EN	<= to_integer(unsigned(h_end));
V_EN	<= to_integer(unsigned(v_end));

--//=======================================================
--//  Structural coding
--//=======================================================

process(v_count,h_count,h_total,h_sync,h_start,h_end,v_total,v_sync,v_start,v_end,v_active_14,v_active_24,v_active_34)
	begin
		h_max 	<= '0';
		hs_end 	<= '0';
		hr_start	<= '0';
		hr_end	<= '0';
		v_max		<= '0';
		vs_end	<= '0';
		vr_start	<= '0';
		vr_end	<= '0';
		v_act_14	<= '0';
		v_act_24	<= '0';
		v_act_34	<= '0';
		if h_count = h_total then h_max <= '1';
		end if;
		if h_count >= h_sync then hs_end <= '1';
		end if;
		if h_count = h_start then hr_start <= '1';
		end if;
		if h_count = h_end then hr_end <= '1';
		end if;
		if v_count = v_total then v_max <= '1';
		end if;
		if v_count >= v_sync then vs_end <= '1';
		end if;
		if v_count = v_start then vr_start <= '1';
		end if;
		if v_count = v_end then vr_end <= '1';
		end if;
		if v_count = v_active_14 then v_act_14 <= '1';
		end if;
		if v_count = v_active_24 then v_act_24 <= '1';  
		end if;
		if v_count = v_active_34 then v_act_34 <= '1';
		end if;
end process;

process (clk,reset_n)
	begin
		if (reset_n='0') then
			Phase <= 0;
		elsif rising_edge(clk) then
			PHASE <= PHASE +1;
			if  PHASE = 1000000 then PHASE <= 0;
			end if;
		end if;
end process;
		

--//horizontal control signals
process (clk,reset_n)
	begin
		if (reset_n='0') then
			h_act_d	<=	'0';
			h_count	<=	(others => '0');
			pixel_x	<=	(others => '0');
			vga_hs	<=	'1';
			h_act		<=	'0';
		elsif rising_edge(clk) then
			h_act_d	<=	h_act;
			if (h_max='1')
				then h_count <=	(others => '0');
				else h_count <=	h_count + "000000000001";
			end if;

			if (h_act_d='1')
				then pixel_x	<=	pixel_x + "00000001";
				else pixel_x	<=	(others => '0');
			end if;
			
			if (PHASE = 0) then PHASE_CNT	<=	PHASE_CNT + "00000001";
			end if;

			if (hs_end='1' and h_max='0')
				then vga_hs	<=	'1';
				else vga_hs	<=	'0';
			end if;
	
			if (hr_start='1')
				then h_act		<=	'1';
				elsif (hr_end='1')
					then h_act	<=	'0';
				end if;
			end if;
	end process;
	

--//vertical control signals
process (clk,reset_n)
	begin
		if (reset_n='0') then
			v_act_d	<=	'0';
			v_count	<=	(others => '0');
			color_mode	<=	(others => '0');
			vga_vs	<=	'1';
			v_act		<=	'0';
		elsif rising_edge(clk) then
			if (h_max='1') then
				v_act_d	  <=	v_act;
				if (v_max='1') then v_count	<=	(others => '0');
									else v_count	<=	v_count + "000000000001";
				end if;
				if (vs_end='1' and v_max='0') then 	vga_vs	<=	'1';
														else	vga_vs	<=	'0';
				end if;
				if (vr_start='1') then	v_act <=	'1';
					elsif (vr_end='1') then	v_act <=	'0';
				end if;
				if (vr_start='1') then color_mode(0) <=	'1';
					elsif (v_act_14='1') then	color_mode(0) <=	'0';
				end if;

				if (v_act_14='1') then	color_mode(1) <=	'1';
					elsif (v_act_24='1') then color_mode(1) <=	'0';
				end if;
				 
				if (v_act_24='1') then	color_mode(2) <=	'1';
					elsif (v_act_34='1') then	color_mode(2) <=	'0';
				end if;
				 
				if (v_act_34='1') then	color_mode(3) <=	'1';
					elsif (vr_end='1') then	color_mode(3) <=	'0';
				end if;
			end if;
		end if;
end process;

--//pattern generator and display enable
process (clk,reset_n)
	begin
		if (reset_n='0') then
			vga_de		<=	'0';
			pre_vga_de	<=	'0';
			boarder		<=	'0';
		elsif rising_edge(clk) then
			vga_de		<=	pre_vga_de;
			pre_vga_de	<=	v_act and h_act;
 
			vga_r <= (others => '0');
			vga_g <= (others => '0');
			vga_b	<= (others => '0');

 
			if ((h_act_d='0' and h_act='1') or hr_end='1' or (v_act_d='0' and v_act='1') or vr_end='1')
				then boarder <='1';
				else boarder <='0';
			end if;
		
			if (boarder='1') then
				vga_r <= (others => '1');
				vga_g <= "00010000";
				vga_b	<= (others => '1');
			end if;

--	display green square if enabled, red if disabled, blue if forced
			for I in 0 to 15 loop
				if ((V_CNT>V_ST+60) and (V_CNT<V_ST+80) and
					(H_CNT>H_ST+150+(20*I)) and (H_CNT<H_ST+150+(20*(I+1)))) then
					if (STATUS(I)='1') then 
						vga_r <= (others => '0');
						vga_g <= (others => '1');
						vga_b	<= (others => '0');
											 else
						vga_r <= (others => '1');
						vga_g <= (others => '0');
						vga_b	<= (others => '0');
					end if;
					if (FORCED(I)='1') then 
						vga_r <= (others => '0');
						vga_g <= (others => '0');
						vga_b	<= (others => '1');
					end if;
				end if;
			end loop;

			
--	display green bar for Power Sourced
				if ((V_CNT>V_ST+120) and (V_CNT<V_ST+140) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+255)) then
						vga_r <= (others => '1');
						vga_g <= (others => '1');
						vga_b	<= (others => '1');
				end if;
				if ((V_CNT>V_ST+120) and (V_CNT<V_ST+140) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+to_integer(unsigned(P_SOURCED)))) then
						vga_r <= (others => '0');
						vga_g <= (others => '1');
						vga_b	<= (others => '0');
				end if;
			

--	display red bar for Power Sinked
				if ((V_CNT>V_ST+150) and (V_CNT<V_ST+170) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+255)) then
						vga_r <= (others => '1');
						vga_g <= (others => '1');
						vga_b	<= (others => '1');
				end if;
				if ((V_CNT>V_ST+150) and (V_CNT<V_ST+170) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+to_integer(unsigned(P_SINKED)))) then
						vga_r <= (others => '1');
						vga_g <= (others => '0');
						vga_b	<= (others => '0');
				end if;

--	display light green bar for Battery Charge
				if ((V_CNT>V_ST+180) and (V_CNT<V_ST+200) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+255)) then
						vga_r <= x"FF";
						vga_g <= (others => '1');
						vga_b	<= (others => '1');
				end if;
				if ((V_CNT>V_ST+180) and (V_CNT<V_ST+200) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+to_integer(unsigned(CHARGE)))) then
						vga_r <= (others => '0');
						vga_g <= x"80";
						vga_b	<= (others => '0');
				end if;

--	display light red bar for Battery Discharge
				if ((V_CNT>V_ST+210) and (V_CNT<V_ST+230) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+255)) then
						vga_r <= x"FF";
						vga_g <= (others => '1');
						vga_b	<= (others => '1');
				end if;
				if ((V_CNT>V_ST+210) and (V_CNT<V_ST+230) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+to_integer(unsigned(DISCHARGE)))) then
						vga_r <= x"80";
						vga_g <= x"00";
						vga_b	<= (others => '0');
				end if;

--	display yellow bar for Battery Status
				if ((V_CNT>V_ST+240) and (V_CNT<V_ST+260) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+255)) then
						vga_r <= x"FF";
						vga_g <= (others => '1');
						vga_b	<= (others => '1');
				end if;
				if ((V_CNT>V_ST+240) and (V_CNT<V_ST+260) and
					(H_CNT>H_ST+180) and (H_CNT<H_ST+180+to_integer(unsigned(BATTERY)))) then
						vga_r <= x"80";
						vga_g <= x"80";
						vga_b	<= x"80";
				end if;

	
--	display logo
				if ((V_CNT>V_ST+300) and (V_CNT<V_ST+420) and
					(H_CNT>H_ST+200) and (H_CNT<H_ST+200+250+1)) then
						if (GIORGI(V_CNT-(V_ST+300+1))(H_CNT-(H_ST+200+1)) = '0') then
							vga_r <= "11111111";--std_logic_vector(to_unsigned(V_CNT-(V_ST+300+1),8));--+PHASE_CNT;
							vga_g <= "11111100"+std_logic_vector(to_unsigned(H_CNT-(H_ST+200+1),8));--+pixel_x;--+PHASE_CNT;
							vga_b	<= "11111000"+ std_logic_vector(to_unsigned(V_CNT-(V_ST+300+1),8))+
										 std_logic_vector(to_unsigned(H_CNT-(H_ST+200+1),8))+PHASE_CNT;
						end if;
				end if;

			
--	display text
				if ((V_CNT>V_ST+120) and (V_CNT<V_ST+136) and
					(H_CNT>H_ST+10) and (H_CNT<H_ST+10+150+1)) then
						if (AVAIL(V_CNT-(V_ST+120+1))(H_CNT-(H_ST+10+1)) = '1') then
							vga_r <= x"ff";
							vga_g <= x"80";
							vga_b	<= x"00";
						end if;
				end if;
		
				if ((V_CNT>V_ST+150) and (V_CNT<V_ST+166) and
					(H_CNT>H_ST+10) and (H_CNT<H_ST+10+150+1)) then
						if (USED(V_CNT-(V_ST+150+1))(H_CNT-(H_ST+10+1)) = '1') then
							vga_r <= x"ff";
							vga_g <= x"80";
							vga_b	<= x"00";
						end if;
				end if;

				if ((V_CNT>V_ST+180) and (V_CNT<V_ST+196) and
					(H_CNT>H_ST+10) and (H_CNT<H_ST+10+150+1)) then
						if (BATCHARGE(V_CNT-(V_ST+180+1))(H_CNT-(H_ST+10+1)) = '1') then
							vga_r <= x"ff";
							vga_g <= x"80";
							vga_b	<= x"00";
						end if;
				end if;

				if ((V_CNT>V_ST+210) and (V_CNT<V_ST+226) and
					(H_CNT>H_ST+10) and (H_CNT<H_ST+10+150+1)) then
						if (BATDISCHARGE(V_CNT-(V_ST+210+1))(H_CNT-(H_ST+10+1)) = '1') then
							vga_r <= x"ff";
							vga_g <= x"80";
							vga_b	<= x"00";
						end if;
				end if;

				if ((V_CNT>V_ST+240) and (V_CNT<V_ST+256) and
					(H_CNT>H_ST+10) and (H_CNT<H_ST+10+150+1)) then
						if (BATSTATUS(V_CNT-(V_ST+240+1))(H_CNT-(H_ST+10+1)) = '1') then
							vga_r <= x"ff";
							vga_g <= x"80";
							vga_b	<= x"00";
						end if;
				end if;

				if ((V_CNT>V_ST+60) and (V_CNT<V_ST+76) and
					(H_CNT>H_ST+10) and (H_CNT<H_ST+10+80+1)) then
						if (LOADS(V_CNT-(V_ST+60+1))(H_CNT-(H_ST+10+1)) = '1') then
							vga_r <= x"ff";
							vga_g <= x"80";
							vga_b	<= x"00";
						end if;
				end if;



--				if ((V_CNT>V_ST+60) and (V_CNT<V_ST+85) and
--					(H_CNT>H_ST+100) and (H_CNT<H_ST+121)) then
--						if (FORNO(((H_CNT-(H_ST+100+1))/8)+V_CNT-(V_ST+60+1))(7-(H_CNT-(H_ST+100+1))+7*((H_CNT-(H_ST+100+1))/8)) ='1') then
--							vga_r <= (others => '1');
--							vga_g <= (others => '1');
--							vga_b	<= (others => '0');
--						end if;
--				end if;




			
--				if (V_CNT>V_ST+30) and (V_CNT<V_ST+50) and
--					(H_CNT>H_ST+100) and (H_CNT<H_ST+120) then
--					vga_r <= (others => '1');
--					vga_g <= (others => '1');
--					vga_b	<= (others => '0');
--				end if;
----
--				if (V_CNT>V_ST+30) and (V_CNT<V_ST+50) and
--					(H_CNT>H_ST+120) and (H_CNT<H_ST+140) then
--					vga_r <= (others => '1');
--					vga_g <= (others => '1');
--					vga_b	<= (others => '0');
--				end if;
--
--				if (V_CNT>V_ST+30) and (V_CNT<V_ST+50) and
--					(H_CNT>H_ST+140) and (H_CNT<H_ST+160) then
--					vga_r <= (others => '1');
--					vga_g <= (others => '1');
--					vga_b	<= (others => '0');
--				end if;
--
--				if (V_CNT>V_ST+30) and (V_CNT<V_ST+50) and
--					(H_CNT>H_ST+100) and (H_CNT<H_ST+120) then
--					vga_r <= (others => '1');
--					vga_g <= (others => '1');
--					vga_b	<= (others => '0');
--				end if;
--
--				if (V_CNT>V_ST+30) and (V_CNT<V_ST+50) and
--					(H_CNT>H_ST+100) and (H_CNT<H_ST+120) then
--					vga_r <= (others => '1');
--					vga_g <= (others => '1');
--					vga_b	<= (others => '0');
--				end if;

					
--			case color_mode is
--				when "0001" =>	vga_r <= pixel_x;
--									vga_g <= (others => '0');
--									vga_b	<= (others => '0');
--									
--				when "0010"	=> vga_g <= pixel_x;
--									vga_r <= (others => '0');
--									vga_b	<= (others => '0');
--									
--				when "0100"	=> vga_b <= pixel_x;
--									vga_g <= (others => '0');
--									vga_r	<= (others => '0');
--									
--				when "1000"	=>	vga_r <= pixel_x;
--									vga_g <= pixel_x;
--									vga_b	<= pixel_x;
--									
--				when others => vga_g <= (others => '0');
--									vga_r <= (others => '0');
--									vga_b <= (others => '0');
--				end case;
	end if;
end process;

end BEH;